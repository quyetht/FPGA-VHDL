LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

entity main is
    port(
        i : in std_logic;
        s : in std_logic_vector(3 downto 0);
        q : out std_
    );