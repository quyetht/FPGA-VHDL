--Viet chuong trinh mo ta VHDL cho mach cong 4 bit khong dau bang cau truc lenh song song
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

entity main is
    port(


    );
end main;

architecture behavi of main is
    begin

    end behavi;
