--viet chuong trinh mo ta VHDL cho mach giai ma nhi phan sang thap phan, sang gray va nguoc lai?

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

entity main is
    port(
        
    );
    end main;

architecture behavi of main is
    begin

    end behavi;