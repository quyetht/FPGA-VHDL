-- viet mo ta VHDL cho IC ghi dich 8 bit hoat dong tai suon duong clock, co tin hieu chot CE muc tich cuc cao
-- tin hieu lap khong dong bo tich cuc cao

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

entity main is
    port(
        

    );
    end main;

architecture behavi of main is
    begin


    end behavi;